library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use STD.ENV.ALL;

entity ALU_TB is
--  Port ( );
end ALU_TB;

architecture Behavioral of ALU_TB is

component ALU is
    port(
        ALUControl : in std_logic_vector(2 downto 0);
        SrcA       : in std_logic_vector(31 downto 0);
        SrcB       : in std_logic_vector(31 downto 0);
        Shamt      : in std_logic_vector(4 downto 0);
        ALUResult  : buffer std_logic_vector(31 downto 0);
        ALUFlags   : out std_logic_vector(3 downto 0)
        );
end component ALU;

signal ALUControl : std_logic_vector(2 downto 0);
signal SrcA       : std_logic_vector(31 downto 0);
signal SrcB       : std_logic_vector(31 downto 0);
signal Shamt      : std_logic_vector(4 downto 0);
signal ALUResult  : std_logic_vector(31 downto 0);
signal ALUFlags   : std_logic_vector(3 downto 0);
        
constant CLK_PERIOD : time := 10 ns;

begin

uut : ALU port map(ALUControl, SrcA, SrcB, Shamt, ALUResult, ALUFlags);

ALUTest : process is
begin
	-- ADD
	ALUControl <= "000"; SrcA <= x"FFFFFFFF"; SrcB <= x"FFFFFFFF"; wait for CLK_PERIOD;
	                     SrcA <= x"00FFFFFF"; SrcB <= x"00ABCD11"; wait for CLK_PERIOD;
						 
	-- SUB
	ALUControl <= "001"; SrcA <= x"FFFFFFFF"; SrcB <= x"FFFFFFFF"; wait for CLK_PERIOD;
	                     SrcA <= x"00FFFFFF"; SrcB <= x"00ABCD11"; wait for CLK_PERIOD;
						 SrcA <= x"FFFFFFFF"; SrcB <= x"0FFFFFFF"; wait for CLK_PERIOD;
			
    -- EOR
	ALUControl <= "010"; SrcA <= x"FFFFFFFF"; SrcB <= x"FFFFFFFF"; wait for CLK_PERIOD;
						 SrcA <= x"00000000"; SrcB <= x"FFFFFFFF"; wait for CLK_PERIOD;
						 SrcA <= x"F0F0F0F0"; SrcB <= x"0F0F0F0F"; wait for CLK_PERIOD;
	
    -- AND	
	ALUControl <= "011"; SrcA <= x"FFFFFFFF"; SrcB <= x"FFFFFFFF"; wait for CLK_PERIOD;
						 SrcA <= x"00000000"; SrcB <= x"FFFFFFFF"; wait for CLK_PERIOD;
						 SrcA <= x"F0F0F0F0"; SrcB <= x"0F0F0F0F"; wait for CLK_PERIOD;
						 
    -- LSL
    ALUControl <= "110"; Shamt <= "00010"; SrcA <= x"0000000F"; wait for CLK_PERIOD;
    
    -- ASR
    ALUControl <= "111"; Shamt <= "00010"; SrcA <= x"0000000F"; wait for CLK_PERIOD;
	
	-- MOV test
	ALUControl <= "100"; SrcB <= x"FFFFFFFF"; wait for CLK_PERIOD;
	
	-- MVN test
	ALUControl <= "101"; wait for CLK_PERIOD;

--	-- CMP test
	ALUControl <= "001"; SrcA <= x"000000F0"; SrcB <= x"0000000F"; wait for CLK_PERIOD;
						 SrcA <= x"0000000F"; SrcB <= x"000000F0"; wait for CLK_PERIOD;
						 SrcA <= x"0000000F"; SrcB <= x"0000000F"; wait for CLK_PERIOD;
						 
	report("Tests completed");
	stop(2);
end process;  
end Behavioral;
